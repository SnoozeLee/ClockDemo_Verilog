module MyClock (
    y,
    x
);
output y;
input x;
Div_100(y, x);
endmodule //MyClock