module Connector (y,x);
output wire y;
input wire x;
assign y = x;
endmodule //Connector